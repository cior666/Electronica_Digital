module AND_compuerta(
    input wire A,
    input wire B,
    output X
);
//logica
assign X=(A & B);
endmodule